library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdram_arbiter_tb is
end sdram_arbiter_tb;

architecture behavior of sdram_arbiter_tb is
begin
end behavior;
